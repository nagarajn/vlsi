////////////////////////////////////////////////////////////////////////////////
// Interface package
////////////////////////////////////////////////////////////////////////////////
//


package intf_pkg;
  `include "intf.sv"
endpackage
