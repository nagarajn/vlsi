////////////////////////////////////////////////////////////////////////////////
// Testbench top level file
////////////////////////////////////////////////////////////////////////////////


//Instantiate the DUT
//Instantiate the VIF
//Instantiate uvm_test

