`define NO_ERR ERR_W'h0

`define ADDR_W 32
`define DATA_W 32

`define ADDR_REG0 `ADDR_W'h0 
`define ADDR_REG1 `ADDR_W'h1 
`define ADDR_REG2 `ADDR_W'h2 
`define ADDR_REG3 `ADDR_W'h3 
`define ADDR_REG4 `ADDR_W'h4 
`define ADDR_REG5 `ADDR_W'h5 
`define ADDR_REG6 `ADDR_W'h6 
`define ADDR_REG7 `ADDR_W'h7 


