`include "intf.sv"
